// Example code for an AHBLite System-on-Chip
//  Iain McNally
//  ECS, University of Soutampton
//
// This module is an AHB-Lite Slave containing one read/write register
//
// Number of addressable locations : 1
// Size of each addressable location : 32 bits
// Supported transfer sizes : Word
// Alignment of base address : Word aligned
//
// Address map :
//   Base addess + 0 : 
//     Read ouput port (oPort) register
//     Write ouput port (oPort) register


`timescale 1ns / 100ps

module ahb_output_port(

  // AHB Global Signals
  input HCLK,
  input HRESETn,

  // AHB Signals from Master to Slave
  input [31:0] HADDR, // With this interface HADDR is ignored
  input [31:0] HWDATA,
  input [2:0] HSIZE,
  input [1:0] HTRANS,
  input HWRITE,
  input HREADY,
  input HSEL,

  // AHB Signals from Slave to Master
  output reg [31:0] HRDATA,
  output HREADYOUT,

  //Non-AHB Signals
  output reg [31:0] oPort

);


  // AHB transfer codes needed in this module
  localparam No_Transfer = 2'b0;

  //control signals are stored in registers
  reg write_enable, read_enable;
 
  //Generate the control signals in the address phase
  always @(posedge HCLK or negedge HRESETn)
    if ( ! HRESETn )
      begin
        write_enable <= 1'b0;
        read_enable <= 1'b0;
      end
    else if ( HREADY && HSEL && (HTRANS != No_Transfer) )
      begin
        write_enable <= HWRITE;
        read_enable <= ! HWRITE;
     end
    else
      begin
        write_enable <= 1'b0;
        read_enable <= 1'b0;
     end

  //Act on control signals in the data phase

  // write
  always @(posedge HCLK or negedge HRESETn)
    if ( ! HRESETn )
      begin
        oPort <= 32'b0;
      end
    else if ( write_enable )
      begin
        oPort <= HWDATA;

        // this is not synthesized but provides useful debugging information
        $display( "oPort: ", HWDATA, " [%x] ", HWDATA, " @", $time );

      end
     
  //read
  always @*
    if ( ! read_enable )
      // (output of zero when not enabled for read is not necessary
      //  but may help with debugging)
      HRDATA = 32'b0;
    else
      HRDATA = oPort;

  //Transfer Response
  assign HREADYOUT = 1'b1; //Single cycle Write & Read. Zero Wait state operations


endmodule

